`timescale 1ns / 1ps

`include "def.v"
module sccomp_dataflow (
    input clk,
    input reset,
    // alu
    output [31:0] a,
    output [31:0] b,
    output [3:0] aluc,
    output [31:0] aluo,
    output zero,
    output carry,
    output negative,
    output overflow,
    // bjudge
    output [31:0] rs,
    output [31:0] rt,
    output [31:0] instr,
    output [31:0] NPC_if_id,
    output B_PC_en,
    output [31:0] B_PC,
    //DMEM
    output [1:0] SC,
    output [2:0] LC,
    output [31:0] Data_in,
    output [31:0] DMEMaddr,
    output CS,
    output DM_W,
    output DM_R,
    input [31:0] Dataout,
    //EX_MEM
    output [3:0] doing_op_id_ex,
    output [31:0] instr_id_ex,
    output [31:0] aluo_ex_mem,
    output [31:0] b_ex_mem,
    output [31:0] instr_ex_mem,
    output [3:0] doing_op_ex_mem,


    //ID_EX
    output [31:0] instr_if_id,
    output [3:0] doing_op ,

    // IF_ID
    output [3:0] jpc_head,
    output [31:0] NPC,
    output [31:0] PC,
    output reg_detect_confict,
    output PC_bobl,
    output JPC_en,
    output [31:0] JPC,
    output halt,

    //IMEM

    //MEM_WB
    output [4:0] rdc,
    output [31:0] rdd,
    output wen ,

    //NPCmaker
    output [31:0] NPC_out,

    //regfile
    output [4:0] rsc,
    output [4:0] rtc,
    output [31:0] rd,
    output [31:0] regfile0,
    output [31:0] regfile1,
    output [31:0] regfile2,
    output [31:0] regfile3,
    output [31:0] regfile4,
    output [31:0] regfile5,
    output [31:0] regfile6,
    output [31:0] regfile7,
    output [31:0] regfile8,
    output [31:0] regfile9,
    output [31:0] regfile10,
    output [31:0] regfile11,
    output [31:0] regfile12,
    output [31:0] regfile13,
    output [31:0] regfile14,
    output [31:0] regfile15,
    output [31:0] regfile16,
    output [31:0] regfile17,
    output [31:0] regfile18,
    output [31:0] regfile19,
    output [31:0] regfile20,
    output [31:0] regfile21,
    output [31:0] regfile22,
    output [31:0] regfile23,
    output [31:0] regfile24,
    output [31:0] regfile25,
    output [31:0] regfile26,
    output [31:0] regfile27,
    output [31:0] regfile28,
    output [31:0] regfile29,
    output [31:0] regfile30,
    output [31:0] regfile31

);
    cpu sccpu(
        .clk(clk),
        .reset(reset),
        .a(a),
        .b(b),
        .aluc(aluc),
        .aluo(aluo),
        .zero(zero),
        .carry(carry),
        .negative(negative),
        .overflow(overflow),
        .rs(rs),
        .rt(rt),
        .instr(instr),
        .NPC_if_id(NPC_if_id),
        .B_PC_en(B_PC_en),
        .B_PC(B_PC),
        .SC(SC),
        .LC(LC),
        .Data_in(Data_in),
        .DMEMaddr(DMEMaddr),
        .CS(CS),
        .DM_W(DM_W),
        .DM_R(DM_R),
        .Dataout(Dataout),
        .doing_op_id_ex(doing_op_id_ex),
        .instr_id_ex(instr_id_ex),
        .aluo_ex_mem(aluo_ex_mem),
        .b_ex_mem(b_ex_mem),
        .instr_ex_mem(instr_ex_mem),
        .doing_op_ex_mem(doing_op_ex_mem),
        .instr_if_id(instr_if_id),
        .doing_op(doing_op),
        .jpc_head(jpc_head),
        .NPC(NPC),
        .PC(PC),
        .reg_detect_confict(reg_detect_confict),
        .PC_bobl(PC_bobl),
        .JPC_en(JPC_en),
        .JPC(JPC),
        .halt(halt),
        .rdc(rdc),
        .rdd(rdd),
        .wen(wen),
        .NPC_out(NPC_out),
        .rsc(rsc),
        .rtc(rtc),
        .rd(rd),
        .regfile0(regfile0),
        .regfile1(regfile1),
        .regfile2(regfile2),
        .regfile3(regfile3),
        .regfile4(regfile4),
        .regfile5(regfile5),
        .regfile6(regfile6),
        .regfile7(regfile7),
        .regfile8(regfile8),
        .regfile9(regfile9),
        .regfile10(regfile10),
        .regfile11(regfile11),
        .regfile12(regfile12),
        .regfile13(regfile13),
        .regfile14(regfile14),
        .regfile15(regfile15),
        .regfile16(regfile16),
        .regfile17(regfile17),
        .regfile18(regfile18),
        .regfile19(regfile19),
        .regfile20(regfile20),
        .regfile21(regfile21),
        .regfile22(regfile22),
        .regfile23(regfile23),
        .regfile24(regfile24),
        .regfile25(regfile25),
        .regfile26(regfile26),
        .regfile27(regfile27),
        .regfile28(regfile28),
        .regfile29(regfile29),
        .regfile30(regfile30),
        .regfile31(regfile31)
    );

    IMEM imem_inst(
        .address(PC),
        .instr_if_id(instr_if_id),
        .instr(instr)
    );

    DMEM dmem_inst(
        .clk(clk),
        .SC(SC),
        .LC(LC),
        .Data_in(Data_in),
        .DMEMaddr(DMEMaddr),
        .CS(CS),
        .DM_W(DM_W),
        .DM_R(DM_R),
        .Dataout(Dataout)
    );

endmodule