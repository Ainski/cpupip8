`include "def.v"
module IMEM(
    input  [31:0] addr,
    output  [31:0] data
);

endmodule